**************************************************************************************
* This is the circuit represneting the spice netlist for nal_nbk_FPGA_ckt_02
*
***************************** written on : Apr 03, 2018 ****************************

r1 1 2 100
r2 1 3 100
r3 2 3 100
r4 2 4 100
r5 3 4 100
i6 3 6 DC 0.002
i7 2 5 DC 0.001
r8 4 5 100
r9 4 6 100
r10 5 6 100
r11 5 7 100
r12 6 7 100
*********************************
r13 3 9 10000 
r14 6 11 10000 
r15 8 9 10000 
r16 8 10 10000 
r17 9 10 10000 
v18 9 11 DC 10
r19 10 12 10000 
r20 11 12 10000 
r21 11 13 10000 
r22 12 13 10000 
r23 10 15 10000
r24 12 17 10000
*****************************8
r25 14 15 100
r26 14 16 100
r27 15 16 100
r28 15 17 100
i29 16 18 DC 0.002
r30 17 18 100
r31 17 19 100
r32 18 19 100
r33 16 20 10000
r34 18 0 10000
v35 20 0 DC 20 
***************************************
.op 
.control
run
print all
.endc

.end

