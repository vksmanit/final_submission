***************************************************************
* NAL_NBK_CKT for FPGA simulation 
***************************************************************
i1 1 2 dc 0.001
r2 1 3 100
r3 2 3 100
r4 2 4 100
r5 3 4 100
*********************************************
r6 3 0 10000
r7 2 5 10000
r8 4 5 10000
r9 4 0 10000
v10 5 0 dc 10
r11 5 6 10000
r12 6 0 10000
**********************************************
.op 
.control
run
print all
.endc

.end

